// vim: set ft=verilog:

`ifndef COLORS_VH_
`define COLORS_VH_

localparam COLOR_BOARD = 12'h985;
localparam COLOR_BG    = 12'h333;
localparam COLOR_BLACK = 12'h111;
localparam COLOR_WHITE = 12'heee;

// magenta-ish color, used to indicate that something's wrong
localparam COLOR_ERROR = 12'he3e;

`endif
